CONFIGURATION cfg OF FILTRO_TD IS
   FOR FILTRO_TEST
      -- default configuration
   END FOR;
END cfg;